-- tb_uart_txd.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_uart_txd is
end tb_uart_txd;

architecture sim of tb_uart_txd is

    -- DUT ��Ʈ�� ����� ��ȣ
    signal rst_l   : std_logic := '0';
    signal clk100m : std_logic := '0';
    signal sw      : std_logic := '0';
    signal txd     : std_logic;

    constant CLK_PERIOD : time := 10 ns;  -- 100MHz (10ns �ֱ�)

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.uart_txd
        port map (
            rst_l   => rst_l,
            clk100m => clk100m,
            sw      => sw,
            txd     => txd
        );

    --------------------------------------------------------------------
    -- 100MHz Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk100m <= '0';
            wait for CLK_PERIOD / 2;
            clk100m <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- ���� + ����ġ �ڱ�
    --------------------------------------------------------------------
    stim_proc : process
    begin
        ----------------------------------------------------------------
        -- 1) �ʱ�: ���� assert (low), ����ġ OFF
        ----------------------------------------------------------------
        rst_l <= '0';
        sw    <= '0';
        wait for 1 us;

        ----------------------------------------------------------------
        -- 2) ���� ����
        ----------------------------------------------------------------
        rst_l <= '1';

        -- PLL lock �� ���� �ʱ�ȭ �ð� ����
        wait for 50 us;

        ----------------------------------------------------------------
        -- 3) ����ġ 1��° Ŭ��
        --    ������ ���� �ð��� ���� ��ư �������� ���� ?s ����
        ----------------------------------------------------------------
        sw <= '1';
        wait for 1 ms;
        sw <= '0';

        -- �� ����('A')�� ���۵� �ð��� ��ٷ� ��
        -- 115200bps���� 1������ �� 87us, �����ְ� 1ms �̻�
        wait for 2 ms;

        ----------------------------------------------------------------
        -- 4) ����ġ 2��° Ŭ��
        ----------------------------------------------------------------
        sw <= '1';
        wait for 1 ms;
        sw <= '0';

        wait for 2 ms;

        ----------------------------------------------------------------
        -- 5) �ùķ��̼� ����
        ----------------------------------------------------------------
        wait;
    end process;

end sim;
