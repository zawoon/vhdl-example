library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SW_INPUT is
    Port (
        rst_l   : in  STD_LOGIC;  -- �ܺ� ���� (Low active)
        clk100m : in  STD_LOGIC;  -- ���� �⺻ 100MHz Ŭ��
        sw      : in  STD_LOGIC;  -- ����ġ �Է�
        led     : out STD_LOGIC   -- LED ���
    );
end SW_INPUT;

architecture Behavioral of SW_INPUT is

    -- Clock Wizard (PLL) ������Ʈ ����
    component my_clk_wiz
        port (
            clk_out1 : out std_logic;
            resetn   : in  std_logic;
            locked   : out std_logic;
            clk_in1  : in  std_logic
        );
    end component;

    signal locked   : std_logic;
    signal clk40m   : std_logic;
    signal rst      : std_logic;

    -- ����ġ ����ȭ �� ��ۿ� ��ȣ
    signal sw_sync1 : std_logic := '0';
    signal sw_sync2 : std_logic := '0';
    signal sw_prev  : std_logic := '0';
    signal led_reg  : std_logic := '0';

begin

    -- 100MHz �� 40MHz Ŭ�� ����
    i_my_clk_wiz : my_clk_wiz
        port map (
            clk_out1 => clk40m,
            resetn   => rst_l,     -- �ܺ� ���� low �� resetn=0
            locked   => locked,
            clk_in1  => clk100m
        );

    -- PLL lock �� �ưų� �ܺ� reset �� ������ rst=1
    rst <= (not locked) or (not rst_l);

    ----------------------------------------------------------------
    -- ����ġ �Է� ����ȭ & ��ư ���� ���� �� LED ���
    ----------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            sw_sync1 <= '0';
            sw_sync2 <= '0';
            sw_prev  <= '0';
            led_reg  <= '0';
        elsif rising_edge(clk40m) then
            -- 2�� ����ȭ(��Ÿ ������ ����)
            sw_sync1 <= sw;
            sw_sync2 <= sw_sync1;

            -- ���� ���¿� ���ؼ� "�տ��� �ڷ�" 0��1 ���ϴ� ���� ����
            if (sw_sync2 = '1') and (sw_prev = '0') then
                led_reg <= not led_reg;   -- ����ġ�� �ѹ� ���� ������ LED ���
            end if;

            -- ���� Ŭ�Ͽ��� ���� ���� �� ����
            sw_prev <= sw_sync2;
        end if;
    end process;

    -- LED ��� ����
    led <= led_reg;

end Behavioral;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SW_INPUT is
    Port (
        rst_l   : in  STD_LOGIC;  -- �ܺ� ���� (Low active)
        clk100m : in  STD_LOGIC;  -- ���� �⺻ 100MHz Ŭ��
        sw      : in  STD_LOGIC;  -- ����ġ �Է�
        led     : out STD_LOGIC   -- LED ���
    );
end SW_INPUT;

architecture Behavioral of SW_INPUT is

    -- Clock Wizard (PLL) ������Ʈ ����
    component my_clk_wiz
        port (
            clk_out1 : out std_logic;
            resetn   : in  std_logic;
            locked   : out std_logic;
            clk_in1  : in  std_logic
        );
    end component;

    signal locked   : std_logic;
    signal clk40m   : std_logic;
    signal rst      : std_logic;

    -- ����ġ ����ȭ �� ��ۿ� ��ȣ
    signal sw_sync1 : std_logic := '0';
    signal sw_sync2 : std_logic := '0';
    signal sw_prev  : std_logic := '0';
    signal led_reg  : std_logic := '0';

begin

    -- 100MHz �� 40MHz Ŭ�� ����
    i_my_clk_wiz : my_clk_wiz
        port map (
            clk_out1 => clk40m,
            resetn   => rst_l,     -- �ܺ� ���� low �� resetn=0
            locked   => locked,
            clk_in1  => clk100m
        );

    -- PLL lock �� �ưų� �ܺ� reset �� ������ rst=1
    rst <= (not locked) or (not rst_l);

    ----------------------------------------------------------------
    -- ����ġ �Է� ����ȭ & ��ư ���� ���� �� LED ���
    ----------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            sw_sync1 <= '0';
            sw_sync2 <= '0';
            sw_prev  <= '0';
            led_reg  <= '0';
        elsif rising_edge(clk40m) then
            -- 2�� ����ȭ(��Ÿ ������ ����)
            sw_sync1 <= sw;
            sw_sync2 <= sw_sync1;

            -- ���� ���¿� ���ؼ� "�տ��� �ڷ�" 0��1 ���ϴ� ���� ����
            if (sw_sync2 = '1') and (sw_prev = '0') then
                led_reg <= not led_reg;   -- ����ġ�� �ѹ� ���� ������ LED ���
            end if;

            -- ���� Ŭ�Ͽ��� ���� ���� �� ����
            sw_prev <= sw_sync2;
        end if;
    end process;

    -- LED ��� ����
    led <= led_reg;

end Behavioral;
