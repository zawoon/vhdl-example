-- SEG7_COUNTER.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SEG7_COUNTER is
    Port (
        rst_l    : in  STD_LOGIC;                  -- �ܺ� ���� (Low active)
        clk100m  : in  STD_LOGIC;                  -- 100MHz �Է� Ŭ��
        sw       : in  STD_LOGIC;                  -- ����ġ �Է�
        seg7     : out STD_LOGIC_VECTOR(6 downto 0) -- a,b,c,d,e,f,g (active-low)
    );
end SEG7_COUNTER;

architecture Behavioral of SEG7_COUNTER is

    --------------------------------------------------------------------
    -- Clock Wizard (PLL) ������Ʈ ����
    --------------------------------------------------------------------
    component my_clk_wiz
        port (
            clk_out1 : out std_logic;  -- ���ο� Ŭ�� (40MHz ��)
            reset    : in  std_logic;  -- Active-high reset
            locked   : out std_logic;  -- PLL lock �÷���
            clk_in1  : in  std_logic   -- 100MHz �Է� Ŭ��
        );
    end component;

    signal locked    : std_logic;
    signal clk40m    : std_logic;                  -- ���� 40MHz Ŭ��
    signal rst       : std_logic;                  -- ���� ���� (High active)

    -- 0~9 ���� ī����
    signal digit_cnt : unsigned(3 downto 0)  := (others => '0');

    signal seg_reg   : std_logic_vector(6 downto 0) := (others => '1');

    -- ����ġ ����ȭ �� edge ����� ��������
    signal sw_sync1  : std_logic := '0';
    signal sw_sync2  : std_logic := '0';
    signal sw_prev   : std_logic := '0';

begin

    --------------------------------------------------------------------
    -- 100MHz �� 40MHz ��ȯ (Clock Wizard �ν��Ͻ�)
    -- reset ��Ʈ�� active-high �̹Ƿ�, low-active�� rst_l�� not �ؼ� ����
    --------------------------------------------------------------------
    i_my_clk_wiz : my_clk_wiz
        port map ( 
            clk_out1 => clk40m,
            reset    => not rst_l,  -- �� �߿�: rst_l�� 1�� �� reset=0 �� �ǵ���
            locked   => locked,
            clk_in1  => clk100m
        );

    -- PLL lock �� �Ǿ��ų�, �ܺ� reset �� ������ rst=1
    rst <= (not locked) or (not rst_l);

    --------------------------------------------------------------------
    -- ����ġ ����(0��1 ��� ����)���� digit_cnt 1 ����
    --------------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            sw_sync1  <= '0';
            sw_sync2  <= '0';
            sw_prev   <= '0';
            digit_cnt <= (others => '0');
        elsif rising_edge(clk40m) then
            -- 2�� ����ȭ (��Ÿ ������ ����)
            sw_sync1 <= sw;
            sw_sync2 <= sw_sync1;

            -- 0��1 ��� ���� ����
            if (sw_sync2 = '1') and (sw_prev = '0') then
                if digit_cnt = 9 then
                    digit_cnt <= (others => '0');
                else
                    digit_cnt <= digit_cnt + 1;
                end if;
            end if;

            -- ���� Ŭ�Ͽ��� ���� ���� ���� ����
            sw_prev <= sw_sync2;
        end if;
    end process;

    --------------------------------------------------------------------
    -- digit_cnt(0~9)�� ���� 7-segment ���� ����
    -- ���� �ֳ��(Common Anode), segment active-low ����
    -- seg7 = "abcdefg"
    --------------------------------------------------------------------
    process(digit_cnt)
    begin
        case digit_cnt is
            when "0000" =>  -- 0
                seg_reg <= "0000001";  -- a,b,c,d,e,f ON, g OFF
            when "0001" =>  -- 1
                seg_reg <= "1001111";  -- b,c ON
            when "0010" =>  -- 2
                seg_reg <= "0010010";
            when "0011" =>  -- 3
                seg_reg <= "0000110";
            when "0100" =>  -- 4
                seg_reg <= "1001100";
            when "0101" =>  -- 5
                seg_reg <= "0100100";
            when "0110" =>  -- 6
                seg_reg <= "0100000";
            when "0111" =>  -- 7
                seg_reg <= "0001111";
            when "1000" =>  -- 8
                seg_reg <= "0000000";
            when "1001" =>  -- 9
                seg_reg <= "0000100";
            when others =>
                seg_reg <= "1111111";  -- blank
        end case;
    end process;

    seg7 <= seg_reg;

end Behavioral;
