-- tb_SEG7_COUNTER_SW.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_SEG7_COUNTER is
end tb_SEG7_COUNTER;

architecture sim of tb_SEG7_COUNTER is

    -- DUT ��Ʈ�� ����� ��ȣ
    signal rst_l   : std_logic := '0';
    signal clk100m : std_logic := '0';
    signal sw      : std_logic := '0';
    signal seg7    : std_logic_vector(6 downto 0);

    constant CLK_PERIOD : time := 10 ns;  -- 100MHz (10ns �ֱ�)

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.SEG7_COUNTER
        port map (
            rst_l   => rst_l,
            clk100m => clk100m,
            sw      => sw,
            seg7    => seg7
        );

    --------------------------------------------------------------------
    -- 100MHz Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk100m <= '0';
            wait for CLK_PERIOD / 2;
            clk100m <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- ���� + ����ġ �ڱ�
    --------------------------------------------------------------------
    stim_proc : process
    begin
        -- �ʱ�: ���� assert (low), ����ġ OFF
        rst_l <= '0';
        sw    <= '0';
        wait for 200 ns;

        -- ���� ����
        rst_l <= '1';

        -- PLL lock �� ���� �ʱ�ȭ �ð� �ణ ��ٸ���
        wait for 2 us;

        ----------------------------------------------------------------
        -- 1��° ��ư Ŭ�� (ª�� �޽�)
        ----------------------------------------------------------------
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        ----------------------------------------------------------------
        -- 2��° Ŭ��
        ----------------------------------------------------------------
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        ----------------------------------------------------------------
        -- 3��° Ŭ��
        ----------------------------------------------------------------
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        ----------------------------------------------------------------
        -- 4��° Ŭ��
        ----------------------------------------------------------------
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        -- �ʿ��ϸ� �� ��������
        -- ...

        -- �ùķ��̼� ����
        wait;
    end process;

end sim;
