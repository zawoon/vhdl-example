library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_spi_master is
end tb_spi_master;

architecture sim of tb_spi_master is

    --------------------------------------------------------------------
    -- DUT�� ����� ��ȣ ����
    --------------------------------------------------------------------
    signal clk       : std_logic := '0';
    signal rst       : std_logic := '1';  -- High active reset

    signal tx_start  : std_logic := '0';
    signal tx_data   : std_logic_vector(7 downto 0) := (others => '0');
    signal tx_busy   : std_logic;

    signal rx_data   : std_logic_vector(7 downto 0);
    signal rx_valid  : std_logic;

    signal sclk      : std_logic;
    signal mosi      : std_logic;
    signal miso      : std_logic := '0';
    signal ss_n      : std_logic;

    --------------------------------------------------------------------
    -- SPI Slave �𵨿� ��ȣ (TB ����)
    --------------------------------------------------------------------
    signal slave_shift : std_logic_vector(7 downto 0) := "10101100";  -- ���� ����

    constant CLK_PERIOD : time := 25 ns;  -- 40MHz �ý��� Ŭ��

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.spi_master
        port map (
            clk      => clk,
            rst      => rst,
            tx_start => tx_start,
            tx_data  => tx_data,
            tx_busy  => tx_busy,
            rx_data  => rx_data,
            rx_valid => rx_valid,
            sclk     => sclk,
            mosi     => mosi,
            miso     => miso,
            ss_n     => ss_n
        );

    --------------------------------------------------------------------
    -- 40MHz �ý��� Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk <= '0';
            wait for CLK_PERIOD/2;
            clk <= '1';
            wait for CLK_PERIOD/2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- ������ SPI Slave ��
    --  - ss_n�� 1 �� idle ����, ���� ������ ���� ���� �ε�
    --  - ss_n�� 0�̰� sclk�� rising edge���� MSB���� �� ��Ʈ�� ����
    --------------------------------------------------------------------
    slave_model : process(sclk, ss_n)
    begin
        if ss_n = '1' then
            -- Slave�� ���� ���·� ���ư��� ���� ���� ���� �ε�
            slave_shift <= "10101100";   -- ���ϴ� ���� (��: 0xAC)
            miso        <= '0';
        elsif rising_edge(sclk) then
            -- MSB���� �� ��Ʈ�� ��������
            miso        <= slave_shift(7);
            slave_shift <= slave_shift(6 downto 0) & '0';
        end if;
    end process;

    --------------------------------------------------------------------
    -- Stimulus ���μ���: ���� ��û �����
    --------------------------------------------------------------------
    stim_proc : process
    begin
        -- 1) �ʱ� ���� Ȱ��
        rst      <= '1';
        tx_start <= '0';
        tx_data  <= (others => '0');
        wait for 1 us;

        -- 2) ���� ����
        rst <= '0';
        wait for 1 us;

        ----------------------------------------------------------------
        -- ù ��° ����: 0x3C ���� ��û
        ----------------------------------------------------------------
        tx_data  <= x"3C";
        tx_start <= '1';
        wait for CLK_PERIOD;
        tx_start <= '0';

        -- ���� �Ϸ���� ��ٸ� (rx_valid�� 1 �Ǵ� �������� ���� ����)
        wait for 500 us;

        ----------------------------------------------------------------
        -- �� ��° ����: 0xA5 ���� ��û
        ----------------------------------------------------------------
        tx_data  <= x"A5";
        tx_start <= '1';
        wait for CLK_PERIOD;
        tx_start <= '0';

        -- �� �� �� �Ϸ� ���
        wait for 500 us;

        -- �ùķ��̼� ����
        wait;
    end process;

end architecture sim;
