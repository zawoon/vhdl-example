library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity spi_master is
    port (
        clk        : in  std_logic;                 -- 40MHz �ý��� Ŭ��
        rst        : in  std_logic;                 -- High active reset

        -- ���� ����
        tx_start   : in  std_logic;                 -- 1 �� ���� ����
        tx_data    : in  std_logic_vector(7 downto 0); -- ������ 8��Ʈ ������
        tx_busy    : out std_logic;                 -- ���� �� = 1

        -- ���� ������
        rx_data    : out std_logic_vector(7 downto 0);
        rx_valid   : out std_logic;

        -- SPI ��ȣ
        sclk       : out std_logic;
        mosi       : out std_logic;
        miso       : in  std_logic;
        ss_n       : out std_logic                  -- Slave Select (active low)
    );
end entity spi_master;

architecture rtl of spi_master is

    --------------------------------------------------------------------
    -- SPI Ŭ�� ���ֱ� (40MHz �� 1MHz)
    -- SCLK_HALF = 20
    -- SCLK = 40MHz / (2 * SCLK_HALF) = 1MHz
    --------------------------------------------------------------------
    constant SCLK_HALF : integer := 20;
    signal div_cnt     : unsigned(7 downto 0) := (others => '0');

    signal sclk_reg  : std_logic := '0';
    signal sclk_div  : std_logic := '0';

    --------------------------------------------------------------------
    -- SPI FSM
    --------------------------------------------------------------------
    type state_t is (IDLE, LOAD, TRANSFER, DONE);
    signal state : state_t := IDLE;

    signal bit_cnt  : unsigned(3 downto 0) := (others => '0');
    signal tx_shift : std_logic_vector(7 downto 0) := (others => '0');
    signal rx_shift : std_logic_vector(7 downto 0) := (others => '0');

begin

    --------------------------------------------------------------------
    -- SCLK ���ֱ� (Mode 0: idle=Low)
    --------------------------------------------------------------------
    process(clk, rst)
    begin
        if rst = '1' then
            div_cnt  <= (others => '0');
            sclk_reg <= '0';
        elsif rising_edge(clk) then
            if state = TRANSFER then
                if div_cnt = SCLK_HALF-1 then
                    div_cnt  <= (others => '0');
                    sclk_reg <= not sclk_reg;    -- toggle SCLK
                else
                    div_cnt <= div_cnt + 1;
                end if;
            else
                sclk_reg <= '0';                 -- IDLE �� Low
                div_cnt  <= (others => '0');
            end if;
        end if;
    end process;

    sclk <= sclk_reg;

    --------------------------------------------------------------------
    -- SPI ���±� (4�ܰ�)
    --------------------------------------------------------------------
    process(clk, rst)
    begin
        if rst = '1' then
            state    <= IDLE;
            ss_n     <= '1';
            tx_busy  <= '0';
            rx_valid <= '0';
            bit_cnt  <= (others => '0');
            tx_shift <= (others => '0');
            rx_shift <= (others => '0');

        elsif rising_edge(clk) then

            rx_valid <= '0';  -- �⺻��

            case state is

                --------------------------------------------------------
                -- 1) IDLE : tx_start�� ��ٸ�
                --------------------------------------------------------
                when IDLE =>
                    ss_n    <= '1';
                    tx_busy <= '0';

                    if tx_start = '1' then
                        state <= LOAD;
                    end if;

                --------------------------------------------------------
                -- 2) LOAD : ���� �غ�
                --------------------------------------------------------
                when LOAD =>
                    ss_n     <= '0';                 -- Slave ����
                    tx_shift <= tx_data;             -- MOSI ����Ʈ �������� �ε�
                    rx_shift <= (others => '0');
                    bit_cnt  <= (others => '0');
                    tx_busy  <= '1';
                    state    <= TRANSFER;

                --------------------------------------------------------
                -- 3) TRANSFER : Mode 0
                --   - SCLK falling edge: MOSI ����
                --   - SCLK rising edge:  MISO ���ø�
                --------------------------------------------------------
                when TRANSFER =>
                    -- Falling edge: MOSI ��� ����
                    if sclk_reg = '0' and div_cnt = 0 then
                        mosi <= tx_shift(7);
                    end if;

                    -- Rising edge: MISO ����
                    if sclk_reg = '1' and div_cnt = 0 then
                        rx_shift <= rx_shift(6 downto 0) & miso;

                        if bit_cnt = 7 then
                            state <= DONE;
                        else
                            bit_cnt <= bit_cnt + 1;
                            tx_shift <= tx_shift(6 downto 0) & '0';
                        end if;
                    end if;

                --------------------------------------------------------
                -- 4) DONE : 1����Ʈ �Ϸ�
                --------------------------------------------------------
                when DONE =>
                    ss_n    <= '1';
                    tx_busy <= '0';
                    rx_valid <= '1';
                    rx_data <= rx_shift;
                    state   <= IDLE;

            end case;
        end if;
    end process;

end architecture rtl;
