library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity uart_txd is
    Port (
        rst_l   : in  STD_LOGIC;   -- �ܺ� ���� (Low active)
        clk100m : in  STD_LOGIC;   -- 100MHz ���� Ŭ��
        sw      : in  STD_LOGIC;   -- ����ġ �Է�
        txd     : out STD_LOGIC    -- UART TX ���
    );
end uart_txd;

architecture Behavioral of uart_txd is

    --------------------------------------------------------------------
    -- Clock Wizard (PLL) ������Ʈ ���� : 100MHz �� 40MHz
    --------------------------------------------------------------------
    component my_clk_wiz
        port (
            clk_out1 : out std_logic;
            resetn   : in  std_logic;
            locked   : out std_logic;
            clk_in1  : in  std_logic
        );
    end component;

    signal clk40m  : std_logic;
    signal locked  : std_logic;
    signal rst     : std_logic;        -- ���� ���� (High active)

    --------------------------------------------------------------------
    -- UART ���� : 115200 bps, 8N1
    -- 40MHz / 115200 �� 347.2  �� ���ְ� 347 ���
    --------------------------------------------------------------------
    constant BAUD_DIV : integer := 347;
    signal baud_cnt   : unsigned(15 downto 0) := (others => '0');
    signal baud_tick  : std_logic := '0';

    --------------------------------------------------------------------
    -- UART �۽� ���±�
    --------------------------------------------------------------------
    type tx_state_t is (IDLE, START_BIT, DATA_BITS, STOP_BIT);
    signal state     : tx_state_t := IDLE;

    signal tx_reg    : std_logic := '1';             -- ���� TX ���� ������ ��
    signal tx_shift  : std_logic_vector(7 downto 0) := (others => '0');
    signal bit_index : unsigned(2 downto 0) := (others => '0');  -- 0~7

    constant TX_DATA_CONST : std_logic_vector(7 downto 0) := x"41";  -- 'A'

    --------------------------------------------------------------------
    -- ����ġ ����ȭ �� ����(����) ����
    --------------------------------------------------------------------
    signal sw_sync1 : std_logic := '0';
    signal sw_sync2 : std_logic := '0';
    signal sw_prev  : std_logic := '0';
    signal sw_pulse : std_logic := '0';  -- 1Ŭ�� �� ��ư �޽�

    --------------------------------------------------------------------
    -- ���� ��û �÷��� (FSM������ ����)
    --------------------------------------------------------------------
    signal tx_req   : std_logic := '0';

begin

    --------------------------------------------------------------------
    -- 100MHz �� 40MHz Ŭ�� ����
    --------------------------------------------------------------------
    i_my_clk_wiz : my_clk_wiz
        port map (
            clk_out1 => clk40m,
            resetn   => rst_l,
            locked   => locked,
            clk_in1  => clk100m
        );

    -- PLL lock �� �Ǿ��ų� �ܺ� reset�� ������ rst=1
    rst <= (not locked) or (not rst_l);

    --------------------------------------------------------------------
    -- ����ġ �Է� ����ȭ + rising edge ���� �� sw_pulse
    --------------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            sw_sync1 <= '0';
            sw_sync2 <= '0';
            sw_prev  <= '0';
            sw_pulse <= '0';
        elsif rising_edge(clk40m) then
            -- 2�� ����ȭ
            sw_sync1 <= sw;
            sw_sync2 <= sw_sync1;

            -- 0 -> 1 ���ϴ� ������ �޽� ����
            if (sw_sync2 = '1') and (sw_prev = '0') then
                sw_pulse <= '1';
            else
                sw_pulse <= '0';
            end if;

            sw_prev <= sw_sync2;
        end if;
    end process;

    --------------------------------------------------------------------
    -- Baud Rate ���ֱ�: 40MHz �� 115200bps (baud_tick ����)
    --------------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            baud_cnt  <= (others => '0');
            baud_tick <= '0';
        elsif rising_edge(clk40m) then
            if baud_cnt = BAUD_DIV - 1 then
                baud_cnt  <= (others => '0');
                baud_tick <= '1';        -- 1 ��Ʈ �Ⱓ���� 1Ŭ�� �޽�
            else
                baud_cnt  <= baud_cnt + 1;
                baud_tick <= '0';
            end if;
        end if;
    end process;

    --------------------------------------------------------------------
    -- UART �۽� ���±� (tx_req�� 1�̸� 1������ ����)
    --------------------------------------------------------------------
    process(clk40m, rst)
    begin
        if rst = '1' then
            state     <= IDLE;
            tx_reg    <= '1';            -- idle �� TX�� High
            tx_shift  <= (others => '0');
            bit_index <= (others => '0');
            tx_req    <= '0';
        elsif rising_edge(clk40m) then

            -- ��ư �޽��� ������ ���� ��û �÷��� �����
            if sw_pulse = '1' then
                tx_req <= '1';
            end if;

            if baud_tick = '1' then
                case state is
                    when IDLE =>
                        tx_reg <= '1';

                        if tx_req = '1' then
                            tx_shift  <= TX_DATA_CONST;       -- 'A' �ε�
                            bit_index <= (others => '0');
                            state     <= START_BIT;
                            tx_req    <= '0';                 -- ��û ����
                        end if;

                    when START_BIT =>
                        -- Start bit: Low
                        tx_reg <= '0';
                        state  <= DATA_BITS;

                    when DATA_BITS =>
                        -- LSB���� 1��Ʈ�� ����
                        tx_reg   <= tx_shift(0);
                        tx_shift <= '0' & tx_shift(7 downto 1);  -- ������ ����Ʈ

                        if bit_index = "111" then   -- 8��Ʈ ���� ��
                            bit_index <= (others => '0');
                            state     <= STOP_BIT;
                        else
                            bit_index <= bit_index + 1;
                        end if;

                    when STOP_BIT =>
                        -- Stop bit: High
                        tx_reg <= '1';
                        state  <= IDLE;

                    when others =>
                        state  <= IDLE;
                        tx_reg <= '1';
                end case;
            end if;
        end if;
    end process;

    --------------------------------------------------------------------
    -- TX ���
    --------------------------------------------------------------------
    txd <= tx_reg;

end Behavioral;

