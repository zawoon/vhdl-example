library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity simple_mcu is
    port (
        clk    : in  std_logic;                          -- �ý��� Ŭ��
        rst_n  : in  std_logic;                          -- active-low reset
        io_out : out std_logic_vector(7 downto 0)        -- LED �� �ܺ� ���
    );
end entity simple_mcu;

architecture rtl of simple_mcu is

    --------------------------------------------------------------------
    -- ROM (Block Memory Generator) ������Ʈ ����
    --------------------------------------------------------------------
    component blk_mem_gen_0
      port (
        clka  : in  std_logic;
        addra : in  std_logic_vector(3 downto 0);
        douta : out std_logic_vector(7 downto 0)
      );
    end component;

    --------------------------------------------------------------------
    -- PC, ALU ������Ʈ ����
    --------------------------------------------------------------------
    component pc_unit
        port (
            clk      : in  std_logic;
            rst_n    : in  std_logic;
            inc_en   : in  std_logic;
            load_en  : in  std_logic;
            load_val  : in  unsigned(3 downto 0);
            pc_out   : out unsigned(3 downto 0)
        );
    end component;

    component alu8
        port (
            acc_in  : in  unsigned(7 downto 0);
            imm     : in  unsigned(7 downto 0);
            opcode  : in  std_logic_vector(3 downto 0);
            acc_out : out unsigned(7 downto 0)
        );
    end component;

    --------------------------------------------------------------------
    -- ���� ����/��ȣ ����
    --------------------------------------------------------------------
    type state_t is (FETCH, EXECUTE);

    signal state   : state_t := FETCH;

    signal pc          : unsigned(3 downto 0) := (others => '0');  -- PC ���
    signal instr       : std_logic_vector(7 downto 0) := (others => '0');
    signal acc         : unsigned(7 downto 0) := (others => '0');  -- ACC
    signal acc_next    : unsigned(7 downto 0) := (others => '0');
    signal out_reg     : std_logic_vector(7 downto 0) := (others => '0');

    -- PC �����
    signal pc_inc_en   : std_logic := '0';
    signal pc_load_en  : std_logic := '0';
    signal pc_load_val : unsigned(3 downto 0) := (others => '0');

begin

    ----------------------------------------------------------------
    -- �ܺ� ���
    ----------------------------------------------------------------
    io_out <= out_reg;

    ----------------------------------------------------------------
    -- Instruction ROM �ν��Ͻ�
    ----------------------------------------------------------------
    u_prog_rom : blk_mem_gen_0
      port map (
        clka  => clk,
        addra => std_logic_vector(pc),
        douta => instr
      );

    ----------------------------------------------------------------
    -- PC �ν��Ͻ�
    ----------------------------------------------------------------
    u_pc : pc_unit
        port map (
            clk      => clk,
            rst_n    => rst_n,
            inc_en   => pc_inc_en,
            load_en  => pc_load_en,
            load_val => pc_load_val,
            pc_out   => pc
        );

    ----------------------------------------------------------------
    -- ALU �ν��Ͻ� (ACC + IMM ���� ����)
    ----------------------------------------------------------------
    -- imm8: 4��Ʈ operand�� 8��Ʈ�� zero-extend
    -- opcode: instr(7 downto 4)
    u_alu : alu8
        port map (
            acc_in  => acc,
            imm     => unsigned("0000" & instr(3 downto 0)),
            opcode  => instr(7 downto 4),
            acc_out => acc_next
        );

    ----------------------------------------------------------------
    -- ������ 2-�������� MCU: FETCH �� EXECUTE
    ----------------------------------------------------------------
    process (clk, rst_n)
        variable opcode  : std_logic_vector(3 downto 0);
        variable operand : std_logic_vector(3 downto 0);
    begin
        if rst_n = '0' then
            state       <= FETCH;
            acc         <= (others => '0');
            out_reg     <= (others => '0');

            pc_inc_en   <= '0';
            pc_load_en  <= '0';
            pc_load_val <= (others => '0');

        elsif rising_edge(clk) then

            -- �⺻��(����Ʈ ����) ����
            pc_inc_en   <= '0';
            pc_load_en  <= '0';
            pc_load_val <= pc_load_val;  -- ����

            case state is

                ----------------------------------------------------
                -- FETCH �ܰ�
                --  - ROM���� instr�� �а�
                --  - PC�� 1 ����
                ----------------------------------------------------
                when FETCH =>
                    pc_inc_en <= '1';     -- �̹� Ŭ�Ͽ� PC <= PC + 1
                    state     <= EXECUTE;

                ----------------------------------------------------
                -- EXECUTE �ܰ�
                ----------------------------------------------------
                when EXECUTE =>
                    opcode  := instr(7 downto 4);
                    operand := instr(3 downto 0);

                    case opcode is

                        when "0000" =>  -- NOP
                            -- ACC ��ȭ ����
                            acc <= acc;  -- (���� ����)

                        when "0001" =>  -- LDI imm : ACC <= imm
                            acc <= acc_next;  -- ALU�� imm �ε�

                        when "0010" =>  -- ADDI imm : ACC <= ACC + imm
                            acc <= acc_next;  -- ALU�� ���� ��� ��ȯ

                        when "0100" =>  -- OUT : out_reg <= ACC
                            out_reg <= std_logic_vector(acc);

                        when "0110" =>  -- JMP addr : PC <= addr
                            pc_load_en  <= '1';
                            pc_load_val <= unsigned(operand);

                        when others =>
                            -- ���ǵ��� ���� opcode �� NOP
                            null;

                    end case;

                    state <= FETCH;

            end case;
        end if;
    end process;

end architecture rtl;

