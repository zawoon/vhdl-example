-- tb_sw_input.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_SW_INPUT is
end tb_SW_INPUT;

architecture sim of tb_SW_INPUT is

    -- DUT ��Ʈ�� ����� ��ȣ��
    signal rst_l   : std_logic := '0';
    signal clk100m : std_logic := '0';
    signal sw      : std_logic := '0';
    signal led     : std_logic;

    constant CLK_PERIOD : time := 10 ns;  -- 100 MHz (10ns �ֱ�)

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.SW_INPUT
        port map (
            rst_l   => rst_l,
            clk100m => clk100m,
            sw      => sw,
            led     => led
        );

    --------------------------------------------------------------------
    -- 100 MHz Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk100m <= '0';
            wait for CLK_PERIOD / 2;
            clk100m <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- ���� + ��ư �Է� �ڱ�
    --------------------------------------------------------------------
    stim_proc : process
    begin
        ----------------------------------------------------------------
        -- �ʱⰪ: ���� assert(��Ȱ��), ����ġ OFF
        ----------------------------------------------------------------
        rst_l <= '0';
        sw    <= '0';
        wait for 200 ns;          -- ���� ����

        ----------------------------------------------------------------
        -- ���� ����
        ----------------------------------------------------------------
        rst_l <= '1';
        -- PLL lock �� �ð� ���� (�뷫 1 us ���� ��ٷ� ��)
        wait for 1 us;

        ----------------------------------------------------------------
        -- ����ġ �Է�: ª�� 0��1��0 �޽��� ���� �� �༭
        -- LED�� ��۵Ǵ��� Ȯ��
        ----------------------------------------------------------------

        -- 1��° Ŭ��
        sw <= '1';
        wait for 200 ns;          -- ��ư ���� �ð�
        sw <= '0';
        wait for 2 us;

        -- 2��° Ŭ��
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        -- 3��° Ŭ��
        sw <= '1';
        wait for 200 ns;
        sw <= '0';
        wait for 2 us;

        -- ���⼭ �ùķ��̼� ����
        wait;
    end process;

end sim;
