library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_simple_mcu is
end tb_simple_mcu;

architecture sim of tb_simple_mcu is

    -- DUT ��Ʈ�� ����� ��ȣ
    signal clk    : std_logic := '0';
    signal rst_n  : std_logic := '0';  -- active-low reset
    signal io_out : std_logic_vector(7 downto 0);

    -- 40MHz �ý��� Ŭ�� (������ 25ns �ֱ�)
    constant CLK_PERIOD : time := 25 ns;

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.simple_mcu
        port map (
            clk    => clk,
            rst_n  => rst_n,
            io_out => io_out
        );

    --------------------------------------------------------------------
    -- 40MHz Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk <= '0';
            wait for CLK_PERIOD / 2;
            clk <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- ���� + ������ ������
    --------------------------------------------------------------------
    stim_proc : process
    begin
        -- ó������ reset assert (rst_n = 0)
        rst_n <= '0';
        wait for 200 ns;

        -- reset ����
        rst_n <= '1';

        -- ����� ���� ������ LED(io_out)�� ����
        -- (Simulation���� ����~���� us ���� ���� ACC�� 1,2,3,... �ö󰡴� �� ����)
        wait for 500 us;

        wait;  -- �ùķ��̼� ����
    end process;

end architecture sim;
