-- tb_uart_rxd.vhd
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_uart_rxd is
end tb_uart_rxd;

architecture sim of tb_uart_rxd is

    --------------------------------------------------------------------
    -- DUT ��Ʈ�� ����� ��ȣ
    --------------------------------------------------------------------
    signal rst_l    : std_logic := '0';
    signal clk100m  : std_logic := '0';
    signal rxd      : std_logic := '1';  -- UART ������ �⺻������ idle=1
    signal rx_data  : std_logic_vector(7 downto 0);
    signal rx_valid : std_logic;

    --------------------------------------------------------------------
    -- Ŭ��/��Ʈ Ÿ�̹� ����
    --------------------------------------------------------------------
    constant CLK100_PERIOD : time := 10 ns;   -- 100MHz
    constant CLK40_PERIOD  : time := 25 ns;   -- 40MHz (Clock Wizard ��� ����)
    constant BAUD_DIV_TB   : integer := 347;  -- ����� ����
    -- 1��Ʈ �Ⱓ (40MHz ���� 347Ŭ��)
    constant BIT_TIME      : time := CLK40_PERIOD * BAUD_DIV_TB;

begin

    --------------------------------------------------------------------
    -- DUT �ν��Ͻ�
    --------------------------------------------------------------------
    uut : entity work.uart_rxd
        port map (
            rst_l    => rst_l,
            clk100m  => clk100m,
            rxd      => rxd,
            rx_data  => rx_data,
            rx_valid => rx_valid
        );

    --------------------------------------------------------------------
    -- 100MHz Ŭ�� ����
    --------------------------------------------------------------------
    clk_gen : process
    begin
        while true loop
            clk100m <= '0';
            wait for CLK100_PERIOD / 2;
            clk100m <= '1';
            wait for CLK100_PERIOD / 2;
        end loop;
    end process;

    --------------------------------------------------------------------
    -- UART �������� ������ִ� ������ procedure
    -- 8N1, LSB first
    --------------------------------------------------------------------
    send_byte_proc : process
        -- �׽�Ʈ�� ���: 'A' = x"41" = 0b0100_0001
        constant TEST_BYTE1 : std_logic_vector(7 downto 0) := x"41"; -- 'A'
        constant TEST_BYTE2 : std_logic_vector(7 downto 0) := x"42"; -- 'B'
    begin
        ----------------------------------------------------------------
        -- 1) �ʱ�: reset assert
        ----------------------------------------------------------------
        rst_l <= '0';
        rxd   <= '1';  -- idle
        wait for 5 us;

        ----------------------------------------------------------------
        -- 2) reset ����
        ----------------------------------------------------------------
        rst_l <= '1';

        -- PLL lock + ���� �ʱ�ȭ ����
        wait for 50 us;

        ----------------------------------------------------------------
        -- 3) ù ��° ����Ʈ ���� : 'A'
        ----------------------------------------------------------------
        -- idle ����
        rxd <= '1';
        wait for BIT_TIME;

        -- Start bit (0)
        rxd <= '0';
        wait for BIT_TIME;

        -- ������ ��Ʈ (LSB first)
        for i in 0 to 7 loop
            rxd <= TEST_BYTE1(i);
            wait for BIT_TIME;
        end loop;

        -- Stop bit (1)
        rxd <= '1';
        wait for BIT_TIME;

        -- ����Ʈ �� ����
        wait for 5 * BIT_TIME;

        ----------------------------------------------------------------
        -- 4) �� ��° ����Ʈ ���� : 'B'
        ----------------------------------------------------------------
        -- Start bit
        rxd <= '0';
        wait for BIT_TIME;

        -- ������ ��Ʈ
        for i in 0 to 7 loop
            rxd <= TEST_BYTE2(i);
            wait for BIT_TIME;
        end loop;

        -- Stop bit
        rxd <= '1';
        wait for BIT_TIME;

        -- ���� idle ����
        wait for 10 * BIT_TIME;

        ----------------------------------------------------------------
        -- 5) �ùķ��̼� ����
        ----------------------------------------------------------------
        wait;
    end process;

end sim;
